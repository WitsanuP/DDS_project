//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.9 Beta-4 Education
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9
//Device Version: C
//Created Time: Sat Jun 22 18:11:50 2024

module coef_prom (dout, clk, oce, ce, reset, ad);

output [47:0] dout;
input clk;
input oce;//Output Clock Enable
input ce; //chip enable
input reset;
input [10:0] ad;

wire [23:0] prom_inst_0_dout_w;
wire [23:0] prom_inst_1_dout_w;
wire [23:0] prom_inst_2_dout_w;
wire [23:0] prom_inst_3_dout_w;
wire [23:0] prom_inst_4_dout_w;
wire [23:0] prom_inst_5_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 8;
defparam prom_inst_0.RESET_MODE = "ASYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h559DDC123E617B8C94938874573101C9873CE78A23B43BB82D98FA53A3EA275B;
defparam prom_inst_0.INIT_RAM_01 = 256'h5CCA2F8BDE27679FCDF10D1F28281F0DF1CC9E6727DD8A2EC95BE363D945A904;
defparam prom_inst_0.INIT_RAM_02 = 256'h9C30BC3EB7268DEA3E89CB043359768A94968E7D634013DD9E5605AA46DA63E4;
defparam prom_inst_0.INIT_RAM_03 = 256'h18D2842CCB61ED71EB5CC42378C40842729AB8CDD9DCD6C6AD8B602CEEA757FE;
defparam prom_inst_0.INIT_RAM_04 = 256'hD0B088561BD78A34D46BF97EF96CD5358CDA1E598BB4D4EBF8FCF7E9D1B18754;
defparam prom_inst_0.INIT_RAM_05 = 256'hC7CDCBBFAA8C6534FBB86C17B951E066E357C1237BCA104C80AACBE3F1F7F3E6;
defparam prom_inst_0.INIT_RAM_06 = 256'hFE2A4E687981807562451FF0B7762BD77A14A42BAA1F8AED4696DD1B507B9EB7;
defparam prom_inst_0.INIT_RAM_07 = 256'h77CA13548AB8DDF80B14140AF8DCB7895212C87519B446CE4EC43195EF4189C8;
defparam prom_inst_0.INIT_RAM_08 = 256'h36AE1D83E0347EC0F8274C697C86877F6E533003CD8D45F39935C751D149B71C;
defparam prom_inst_0.INIT_RAM_09 = 256'h3CDA6FFA7DF667CE2B80CC0E47779EBBD0DBDDD6C6AC895E29EAA352F9962AB4;
defparam prom_inst_0.INIT_RAM_0A = 256'h8B4F0ABB63029825A82394FC5BB0FD407AABD3F10713161001E8C69C682AE494;
defparam prom_inst_0.INIT_RAM_0B = 256'h2711F1C8965A16C87111A835BA35A71070C6135893C5ED0D2330342F2109E8BE;
defparam prom_inst_0.INIT_RAM_0C = 256'h132227241701E2BA894E0ABD6708A02EB32FA20C6CC4125793C5EF0F26343935;
defparam prom_inst_0.INIT_RAM_0D = 256'h5186B0D2EBFA01FEF2DDBE97662CE99D48E98111971387F153ABFA407CB0DAFB;
defparam prom_inst_0.INIT_RAM_0E = 256'hE63F8FD614497597B0C0C7C5BAA5876130F7B56915B750E066E458C3257ECE14;
defparam prom_inst_0.INIT_RAM_0F = 256'hD351C73396F04189C7FC284B65767D7C715D4019EAB16F24D0730D9D24A21783;
defparam prom_inst_0.INIT_RAM_10 = 256'h1DC15BED75F46AD63A94E52D6CA2CFF20C1D25241A06E9C4955C1BD17D20BA4B;
defparam prom_inst_0.INIT_RAM_11 = 256'hC8915006B357F2840C8B026FD22D7FC7063C698DA8B9C2C1B7A4876233FBBB70;
defparam prom_inst_0.INIT_RAM_12 = 256'hD8C5A984561FDE9542E681139C1B92FF63BE105898CEFB1F3A4C55544A381CF6;
defparam prom_inst_0.INIT_RAM_13 = 256'h50626A6A614E320EDFA8681FCC700B9D26A61C8AEE499BE4245A87ACC7D9E1E1;
defparam prom_inst_0.INIT_RAM_14 = 256'h346B98BDD8EAF3F2E9D6BA966830F0A754F89426AE2EA51276D2246CACE31034;
defparam prom_inst_0.INIT_RAM_15 = 256'h8BE53780BFF6234762747D7C7360441FF1BA7930DD811CAE37B72D9BFF5AACF5;
defparam prom_inst_0.INIT_RAM_16 = 256'h57D64CB91C77C9115086B3D7F2040C0B02EFD3AD7F4807BD6A0EA93BC443B926;
defparam prom_inst_0.INIT_RAM_17 = 256'h9D40DA6BF372E854B81263ABEA204C708A9BA3A29885694314DD9C52FFA23DCE;
defparam prom_inst_0.INIT_RAM_18 = 256'h632AE89D49EC85169D1C91FD60B90A5190C5F1142E3F46453A270AE4B57C3BF1;
defparam prom_inst_0.INIT_RAM_19 = 256'hAE987A5323E9A75B06A841D158D54AB51770C007457AA5C8E1F1F8F6EBD7B993;
defparam prom_inst_0.INIT_RAM_1A = 256'h8290969286705129F7BD7A2DD87911A026A31781E33B8AD00D416C8EA6B6BCB9;
defparam prom_inst_0.INIT_RAM_1B = 256'hE51740607784898477604017E5AA6518C162F9870C88FB64C51C6BB0EC1F496A;
defparam prom_inst_0.INIT_RAM_1C = 256'hDD337FC2FC2D557389959993846D4C21EEB26D1EC666FC890D88FA62C21866AA;
defparam prom_inst_0.INIT_RAM_1D = 256'h70E857BE1B6FBAFC34648BA8BCC8CAC3B39A784C18DA9444EB891EAA2DA7177F;
defparam prom_inst_0.INIT_RAM_1E = 256'hA33ED059D950BE237FD11B5B92C1E602151F1F1706EBC89B6526DE8D33D064EE;
defparam prom_inst_0.INIT_RAM_1F = 256'h7C3AEF9A3DD768EF6DE34FB20C5DA5E41A476A85969F9E9481654012DA9A51FE;
defparam prom_inst_0.INIT_RAM_20 = 256'h01E2B9884D09BC66079F2EB431A40F70C9185E9BCFFA1C35454B493D290BE4B5;
defparam prom_inst_0.INIT_RAM_21 = 256'h3A3D37270FEDC38F530DBE66059B28AC27990161B7054984B7E0001725292518;
defparam prom_inst_0.INIT_RAM_22 = 256'h2C516D80898A8270563206D09149F89E3BCF5ADC55C42B88DD286BA4D4FB192E;
defparam prom_inst_0.INIT_RAM_23 = 256'hDE256398C3E6FF1017160BF7DBB5864E0DC37013AE40C848BE2C90EB3E87C7FE;
defparam prom_inst_0.INIT_RAM_24 = 256'h58C02076C30843759EBED5E3E8E4D7C1A279480ECA7E28C962F177F468D4368E;
defparam prom_inst_0.INIT_RAM_25 = 256'h9F29AA2290F653A7F1336C9BC2DFF3FF01FAEAD2B0855114CE7F27C55BE86BE6;
defparam prom_inst_0.INIT_RAM_26 = 256'hBB6709A232B937AC187BD5256DACE20E324D5E67665D4A2E0ADCA5651DCB700C;
defparam prom_inst_0.INIT_RAM_27 = 256'hB48144FEAF57F68C199D188AF353A9F73C78AAD4F40C1B201D10FBDCB4844A07;
defparam prom_inst_0.INIT_RAM_28 = 256'h927E623D0FD8984FFCA13DD059DA52C02683D621629BCAF10E222E30291A01DF;
defparam prom_inst_0.INIT_RAM_29 = 256'h5A686C685A4424FBCA8F4BFFA94AE372F875E955B71060A7E51A476A84959D9C;
defparam prom_inst_0.INIT_RAM_2A = 256'h1745698598A1A29A896E4B1FE9AB6413BA57EC78FA74E44CAA004D90CBFC2544;
defparam prom_inst_0.INIT_RAM_2B = 256'hCF1D619DD0FA1A32414743372204DDAC7331E69134CE5FE665DB48AB0658A1E0;
defparam prom_inst_0.INIT_RAM_2C = 256'h8BF85DB80B5495CDFB213D515B5D56452C0ADEAA6D26D77F1DB340C33EB01978;
defparam prom_inst_0.INIT_RAM_2D = 256'h53E064DF51BA1A71BF0440749EBFD7E6EDEADECAAC85561DDB913DE17B0C9514;
defparam prom_inst_0.INIT_RAM_2E = 256'h2FDB7F19AA32B22896FA56A8F2326A98BEDAEEF9FBF3E3CAA87C480BC5761EBD;
defparam prom_inst_0.INIT_RAM_2F = 256'h29F4B66F20C765FB870B85F75FBF1563A8E316406179888E8A7E694B25F5BC7A;
defparam prom_inst_0.INIT_RAM_30 = 256'h483213EBBA803DF19C3FD868EF6EE350B30E5FA8E81E4C718DA0AAAAA2917855;
defparam prom_inst_0.INIT_RAM_31 = 256'h979F9E9582674215DE9F5706AB48DC67E962D23A98ED397DB7E9113147555A56;
defparam prom_inst_0.INIT_RAM_32 = 256'h1E44617681847E6E56350BD89C5709B253EA78FE7AEE59BA1363AAE81C496C86;
defparam prom_inst_0.INIT_RAM_33 = 256'hE62A6597C1E1F9070D0AFDE8CAA3733BF9AE5AFE982AB332A9177CD82B75B6EE;
defparam prom_inst_0.INIT_RAM_34 = 256'hF85AB3034A88BDE90C26384040372409E5B88243FBAB51EE830E910B7CE34298;
defparam prom_inst_0.INIT_RAM_35 = 256'h60DF54C22681D31D5D95C4E9061A25282111F9D7AD793DF8AA53F38A189E1A8E;
defparam prom_inst_0.INIT_RAM_36 = 256'h25C154DE5FD746AD0A5FABED275880A0B6C3C8C3B6A0815928EEAB5F0BAD47D8;
defparam prom_inst_0.INIT_RAM_37 = 256'h530BBA61FF9420A31D8EF756ADFA3F7BAED8FA122128261A06E9C3955D1CD380;
defparam prom_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000474F4F463318F4C791;
defparam prom_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[23:0],dout[15:8]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 8;
defparam prom_inst_1.RESET_MODE = "ASYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h4149515A626A727A828A929AA2AAB2B9C1C9D0D8E0E7EFF6FE050C141B222A31;
defparam prom_inst_1.INIT_RAM_01 = 256'h252E38414A545D666F78828B949DA6AFB7C0C9D2DBE3ECF5FD060E171F283039;
defparam prom_inst_1.INIT_RAM_02 = 256'hE4EFF9040E19232D38424C57616B757F89939DA7B1BBC5CED8E2ECF5FF08121B;
defparam prom_inst_1.INIT_RAM_03 = 256'h7F8A96A2ADB9C4D0DBE7F2FE0914202B36414C57626D78838E99A4AFB9C4CFD9;
defparam prom_inst_1.INIT_RAM_04 = 256'hF4010E1B2834414E5A6773808C99A5B2BECAD7E3EFFB07131F2B37434F5B6773;
defparam prom_inst_1.INIT_RAM_05 = 256'h4553616F7D8B99A7B4C2D0DEEBF90614212F3C4A5764727F8C99A6B3C0CDDAE7;
defparam prom_inst_1.INIT_RAM_06 = 256'h7181909FAEBDCCDBEAF9081625344351606F7D8C9AA9B7C5D4E2F0FF0D1B2937;
defparam prom_inst_1.INIT_RAM_07 = 256'h79899AAABACADAEAFB0B1B2B3A4A5A6A7A8A99A9B9C8D8E7F706162534445362;
defparam prom_inst_1.INIT_RAM_08 = 256'h5C6D7F90A1B3C4D5E6F8091A2B3C4D5E6F8091A2B2C3D4E4F506162737485869;
defparam prom_inst_1.INIT_RAM_09 = 256'h1A2C3F516476899BAEC0D2E5F7091B2D3F5163758799ABBDCFE0F2041527394A;
defparam prom_inst_1.INIT_RAM_0A = 256'hB3C7DBEE0216293D5064778A9EB1C4D8EBFE1124384B5E718496A9BCCFE2F407;
defparam prom_inst_1.INIT_RAM_0B = 256'h283D51667B90A5B9CEE3F70C2035495E72869BAFC3D7EB0014283C5064788B9F;
defparam prom_inst_1.INIT_RAM_0C = 256'h788EA4BAD0E6FB11273D53687E94A9BFD4EAFF152A3F556A7F94A9BFD4E9FE13;
defparam prom_inst_1.INIT_RAM_0D = 256'hA3BAD1E8FF162E445B7289A0B7CEE4FB12283F566C8399AFC6DCF2091F354B61;
defparam prom_inst_1.INIT_RAM_0E = 256'hA9C2DAF20B233B536B839BB3CBE3FB132B425A728AA1B9D0E8FF172E465D748C;
defparam prom_inst_1.INIT_RAM_0F = 256'h8BA5BED8F10A243D566F89A2BBD4ED061F38516A829BB4CDE5FE172F48607991;
defparam prom_inst_1.INIT_RAM_10 = 256'h49637E98B3CDE8021D37516C86A0BAD4EF09233D57718AA4BED8F20B253F5872;
defparam prom_inst_1.INIT_RAM_11 = 256'hE1FD1935506C87A3BFDAF6112C48637E9AB5D0EB06213C57728DA8C3DEF8132E;
defparam prom_inst_1.INIT_RAM_12 = 256'h55728FACC9E6021F3C587592AECBE703203C597591ADC9E6021E3A56728EAAC5;
defparam prom_inst_1.INIT_RAM_13 = 256'hA5C3E1FF1D3B597794B2D0EE0B294764829FBDDAF715324F6D8AA7C4E1FE1B38;
defparam prom_inst_1.INIT_RAM_14 = 256'hD0EF0E2D4C6B8AA9C8E70625446381A0BFDDFC1B39587695B3D1F00E2C4A6987;
defparam prom_inst_1.INIT_RAM_15 = 256'hD6F61737577798B8D8F81838587898B8D7F71737567696B5D5F41433527291B0;
defparam prom_inst_1.INIT_RAM_16 = 256'hB8D9FB1C3E5F80A2C3E4052647698AABCCEC0D2E4F7091B1D2F31334547595B6;
defparam prom_inst_1.INIT_RAM_17 = 256'h7598BADDFF22446789ACCEF0123557799BBDDF0123456789ABCCEE1031537596;
defparam prom_inst_1.INIT_RAM_18 = 256'h0E3255799DC0E4082B4F7295B9DC002346698CB0D3F6193C5F82A5C7EA0D3052;
defparam prom_inst_1.INIT_RAM_19 = 256'h82A7CCF1163A5F84A9CDF2163B5F84A8CDF1153A5E82A6CAEE12365A7EA2C6EA;
defparam prom_inst_1.INIT_RAM_1A = 256'hD2F81E446A90B6DC01274D7398BEE4092F547A9FC4EA0F345A7FA4C9EE13385D;
defparam prom_inst_1.INIT_RAM_1B = 256'hFD254C739AC1E80F365D84ABD1F81F466C93B9E0072D537AA0C7ED13396086AC;
defparam prom_inst_1.INIT_RAM_1C = 256'h042D557DA5CEF61E466E96BEE60E365E85ADD5FD244C739BC3EA11396088AFD6;
defparam prom_inst_1.INIT_RAM_1D = 256'hE7103A638DB6DF08325B84ADD6FF28517AA3CCF51E466F98C0E9123A638BB4DC;
defparam prom_inst_1.INIT_RAM_1E = 256'hA5D0FA254F7AA4CFF9234E78A2CCF6214B759FC9F31C46709AC4ED17416A94BD;
defparam prom_inst_1.INIT_RAM_1F = 256'h3F6B96C2EE1945709CC7F31E4A75A0CBF7224D78A3CEF9244F7AA5D0FA25507A;
defparam prom_inst_1.INIT_RAM_20 = 256'hB5E10E3B6895C1EE1B4774A0CDF926527EABD7032F5B88B4E00C386490BCE713;
defparam prom_inst_1.INIT_RAM_21 = 256'h06346290BEEB194775A3D0FE2C5987B4E20F3D6A97C5F21F4C79A7D4012E5B88;
defparam prom_inst_1.INIT_RAM_22 = 256'h336291C0EF1E4D7CABDA09376695C3F2214F7EACDB09386694C3F11F4D7BAAD8;
defparam prom_inst_1.INIT_RAM_23 = 256'h3B6C9CCCFC2C5C8DBDED1D4C7CACDC0C3C6B9BCBFA2A5989B8E8174676A5D403;
defparam prom_inst_1.INIT_RAM_24 = 256'h205183B4E5174879AADB0C3D6E9FD001326394C5F5265787B8E819497AAADB0B;
defparam prom_inst_1.INIT_RAM_25 = 256'hE0134578AADC0F4173A6D80A3C6EA0D20536689ACCFE306293C5F7285A8BBDEE;
defparam prom_inst_1.INIT_RAM_26 = 256'h7CB0E4174B7EB2E5194C7FB3E6194C80B3E6194C7FB2E5184B7DB0E316487BAE;
defparam prom_inst_1.INIT_RAM_27 = 256'hF4295E92C7FC30659ACE03376BA0D4083D71A5D90D4276AADE124579ADE11549;
defparam prom_inst_1.INIT_RAM_28 = 256'h487EB4EA20558BC1F62C6297CD02386DA3D80D4378ADE2174D82B7EC21568BBF;
defparam prom_inst_1.INIT_RAM_29 = 256'h78AFE61D548BC2F82F669DD30A4177AEE41B5188BEF52B6197CE043A70A6DC12;
defparam prom_inst_1.INIT_RAM_2A = 256'h84BCF42C649CD40C447CB4EC235B93CB023A71A9E0184F87BEF62D649BD20A41;
defparam prom_inst_1.INIT_RAM_2B = 256'h6BA5DE175089C3FC356EA7E019528AC3FC356DA6DF175088C1F9326AA3DB134B;
defparam prom_inst_1.INIT_RAM_2C = 256'h2F69A4DE19538DC7013C76B0EA245E98D20C457FB9F32C66A0D9134C86BFF932;
defparam prom_inst_1.INIT_RAM_2D = 256'hCF0A4681BDF8346FAAE6215C97D20D4883BEF9346FAAE5205A95D00A4580BAF5;
defparam prom_inst_1.INIT_RAM_2E = 256'h4B87C4013D7AB6F32F6BA8E4205D99D5114D89C5013D79B5F12D69A5E01C5893;
defparam prom_inst_1.INIT_RAM_2F = 256'hA3E01E5C9AD7155290CE0B4886C3013E7BB8F63370ADEA2764A1DE1B5894D10E;
defparam prom_inst_1.INIT_RAM_30 = 256'hD7165593D211508ECD0C4A89C7064483C1003E7CBAF93775B3F12F6DABE92765;
defparam prom_inst_1.INIT_RAM_31 = 256'hE72767A7E72767A7E62666A6E52564A4E32362A2E120609FDE1D5D9CDB1A5998;
defparam prom_inst_1.INIT_RAM_32 = 256'hD4155697D8195A9BDC1D5E9EDF2061A1E22263A3E42465A5E62666A6E72767A7;
defparam prom_inst_1.INIT_RAM_33 = 256'h9CDF2163A5E7296CAEF03173B5F7397BBCFE4081C3054688C90B4C8DCF105192;
defparam prom_inst_1.INIT_RAM_34 = 256'h4185C80C4F92D5185C9FE22568ABEE3173B6F93C7EC1044689CC0E5193D5185A;
defparam prom_inst_1.INIT_RAM_35 = 256'hC3074C90D5195DA2E62A6EB2F73B7FC3074B8ED2165A9EE12569ACF03477BBFE;
defparam prom_inst_1.INIT_RAM_36 = 256'h2166ACF1377CC2074D92D71C62A7EC3176BB00458ACF14599EE2276CB1F53A7E;
defparam prom_inst_1.INIT_RAM_37 = 256'h5BA2E82F75BC034990D61C63A9EF367CC2084E95DB2167ADF3387EC40A5095DB;
defparam prom_inst_1.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000DD246BB2F94086CD14;
defparam prom_inst_1.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[23:0],dout[23:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 8;
defparam prom_inst_2.RESET_MODE = "ASYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'hFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFDFDFDFDFDFDFD;
defparam prom_inst_2.INIT_RAM_01 = 256'hFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFCFCFCFCFCFCFC;
defparam prom_inst_2.INIT_RAM_02 = 256'hF9F9F9FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFBFBFB;
defparam prom_inst_2.INIT_RAM_03 = 256'hF8F8F8F8F8F8F8F8F8F8F8F8F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9;
defparam prom_inst_2.INIT_RAM_04 = 256'hF6F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F8F8F8F8F8F8F8F8F8F8;
defparam prom_inst_2.INIT_RAM_05 = 256'hF5F5F5F5F5F5F5F5F5F5F5F5F5F5F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6;
defparam prom_inst_2.INIT_RAM_06 = 256'hF3F3F3F3F3F3F3F3F3F3F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F5F5F5F5;
defparam prom_inst_2.INIT_RAM_07 = 256'hF1F1F1F1F1F1F1F1F1F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F3F3F3F3F3F3F3;
defparam prom_inst_2.INIT_RAM_08 = 256'hEFEFEFEFEFEFEFEFEFEFF0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F1F1F1F1F1F1F1;
defparam prom_inst_2.INIT_RAM_09 = 256'hEDEDEDEDEDEDEDEDEDEDEDEDEDEEEEEEEEEEEEEEEEEEEEEEEEEEEEEFEFEFEFEF;
defparam prom_inst_2.INIT_RAM_0A = 256'hEAEAEAEAEBEBEBEBEBEBEBEBEBEBEBEBEBEBECECECECECECECECECECECECECED;
defparam prom_inst_2.INIT_RAM_0B = 256'hE8E8E8E8E8E8E8E8E8E8E8E9E9E9E9E9E9E9E9E9E9E9E9EAEAEAEAEAEAEAEAEA;
defparam prom_inst_2.INIT_RAM_0C = 256'hE5E5E5E5E5E5E5E6E6E6E6E6E6E6E6E6E6E6E6E7E7E7E7E7E7E7E7E7E7E7E7E8;
defparam prom_inst_2.INIT_RAM_0D = 256'hE2E2E2E2E2E3E3E3E3E3E3E3E3E3E3E3E4E4E4E4E4E4E4E4E4E4E4E5E5E5E5E5;
defparam prom_inst_2.INIT_RAM_0E = 256'hDFDFDFDFE0E0E0E0E0E0E0E0E0E0E0E1E1E1E1E1E1E1E1E1E1E1E2E2E2E2E2E2;
defparam prom_inst_2.INIT_RAM_0F = 256'hDCDCDCDCDCDDDDDDDDDDDDDDDDDDDDDEDEDEDEDEDEDEDEDEDEDEDFDFDFDFDFDF;
defparam prom_inst_2.INIT_RAM_10 = 256'hD9D9D9D9D9D9D9DADADADADADADADADADADBDBDBDBDBDBDBDBDBDBDCDCDCDCDC;
defparam prom_inst_2.INIT_RAM_11 = 256'hD5D5D6D6D6D6D6D6D6D6D6D7D7D7D7D7D7D7D7D7D8D8D8D8D8D8D8D8D8D8D9D9;
defparam prom_inst_2.INIT_RAM_12 = 256'hD2D2D2D2D2D2D3D3D3D3D3D3D3D3D3D4D4D4D4D4D4D4D4D4D5D5D5D5D5D5D5D5;
defparam prom_inst_2.INIT_RAM_13 = 256'hCECECECECFCFCFCFCFCFCFCFD0D0D0D0D0D0D0D0D0D1D1D1D1D1D1D1D1D1D2D2;
defparam prom_inst_2.INIT_RAM_14 = 256'hCACACBCBCBCBCBCBCBCBCCCCCCCCCCCCCCCCCCCDCDCDCDCDCDCDCDCECECECECE;
defparam prom_inst_2.INIT_RAM_15 = 256'hC6C6C7C7C7C7C7C7C7C7C8C8C8C8C8C8C8C8C9C9C9C9C9C9C9C9CACACACACACA;
defparam prom_inst_2.INIT_RAM_16 = 256'hC2C2C2C3C3C3C3C3C3C3C4C4C4C4C4C4C4C4C5C5C5C5C5C5C5C5C6C6C6C6C6C6;
defparam prom_inst_2.INIT_RAM_17 = 256'hBEBEBEBEBEBFBFBFBFBFBFBFC0C0C0C0C0C0C0C1C1C1C1C1C1C1C1C2C2C2C2C2;
defparam prom_inst_2.INIT_RAM_18 = 256'hBABABABABABABABBBBBBBBBBBBBBBCBCBCBCBCBCBCBCBDBDBDBDBDBDBDBEBEBE;
defparam prom_inst_2.INIT_RAM_19 = 256'hB5B5B5B5B6B6B6B6B6B6B6B7B7B7B7B7B7B7B8B8B8B8B8B8B8B9B9B9B9B9B9B9;
defparam prom_inst_2.INIT_RAM_1A = 256'hB0B0B1B1B1B1B1B1B2B2B2B2B2B2B2B3B3B3B3B3B3B3B4B4B4B4B4B4B4B5B5B5;
defparam prom_inst_2.INIT_RAM_1B = 256'hABACACACACACACADADADADADADADAEAEAEAEAEAEAFAFAFAFAFAFAFB0B0B0B0B0;
defparam prom_inst_2.INIT_RAM_1C = 256'hA7A7A7A7A7A7A7A8A8A8A8A8A8A9A9A9A9A9A9A9AAAAAAAAAAAAABABABABABAB;
defparam prom_inst_2.INIT_RAM_1D = 256'hA1A2A2A2A2A2A2A3A3A3A3A3A3A3A4A4A4A4A4A4A5A5A5A5A5A5A6A6A6A6A6A6;
defparam prom_inst_2.INIT_RAM_1E = 256'h9C9C9C9D9D9D9D9D9D9E9E9E9E9E9E9F9F9F9F9F9FA0A0A0A0A0A0A1A1A1A1A1;
defparam prom_inst_2.INIT_RAM_1F = 256'h97979797979898989898989999999999999A9A9A9A9A9A9B9B9B9B9B9B9C9C9C;
defparam prom_inst_2.INIT_RAM_20 = 256'h9191929292929292939393939393949494949495959595959596969696969697;
defparam prom_inst_2.INIT_RAM_21 = 256'h8C8C8C8C8C8C8D8D8D8D8D8D8E8E8E8E8E8F8F8F8F8F8F909090909091919191;
defparam prom_inst_2.INIT_RAM_22 = 256'h8686868686878787878788888888888889898989898A8A8A8A8A8A8B8B8B8B8B;
defparam prom_inst_2.INIT_RAM_23 = 256'h8080808080818181818182828282828383838383838484848484858585858586;
defparam prom_inst_2.INIT_RAM_24 = 256'h7A7A7A7A7A7B7B7B7B7B7C7C7C7C7C7D7D7D7D7D7D7E7E7E7E7E7F7F7F7F7F80;
defparam prom_inst_2.INIT_RAM_25 = 256'h7374747474747575757575767676767677777777777778787878787979797979;
defparam prom_inst_2.INIT_RAM_26 = 256'h6D6D6D6E6E6E6E6E6F6F6F6F6F70707070707171717171727272727273737373;
defparam prom_inst_2.INIT_RAM_27 = 256'h6667676767676868686869696969696A6A6A6A6A6B6B6B6B6B6C6C6C6C6C6D6D;
defparam prom_inst_2.INIT_RAM_28 = 256'h6060606061616161616262626263636363636464646464656565656566666666;
defparam prom_inst_2.INIT_RAM_29 = 256'h5959595A5A5A5A5A5B5B5B5B5C5C5C5C5C5D5D5D5D5D5E5E5E5E5F5F5F5F5F60;
defparam prom_inst_2.INIT_RAM_2A = 256'h5252525353535354545454545555555556565656565757575757585858585959;
defparam prom_inst_2.INIT_RAM_2B = 256'h4B4B4B4C4C4C4C4C4D4D4D4D4E4E4E4E4E4F4F4F4F5050505050515151515252;
defparam prom_inst_2.INIT_RAM_2C = 256'h44444444454545454646464646474747474848484848494949494A4A4A4A4A4B;
defparam prom_inst_2.INIT_RAM_2D = 256'h3C3D3D3D3D3D3E3E3E3E3F3F3F3F404040404041414141424242424343434343;
defparam prom_inst_2.INIT_RAM_2E = 256'h35353536363636363737373738383838393939393A3A3A3A3A3B3B3B3B3C3C3C;
defparam prom_inst_2.INIT_RAM_2F = 256'h2D2D2E2E2E2E2F2F2F2F30303030313131313132323232333333333434343435;
defparam prom_inst_2.INIT_RAM_30 = 256'h25262626262727272728282828292929292A2A2A2A2A2B2B2B2B2C2C2C2C2D2D;
defparam prom_inst_2.INIT_RAM_31 = 256'h1D1E1E1E1E1F1F1F1F2020202021212121222222222323232324242424252525;
defparam prom_inst_2.INIT_RAM_32 = 256'h15161616161717171718181818191919191A1A1A1A1B1B1B1B1C1C1C1C1D1D1D;
defparam prom_inst_2.INIT_RAM_33 = 256'h0D0D0E0E0E0E0F0F0F0F10101010111111111212121313131314141414151515;
defparam prom_inst_2.INIT_RAM_34 = 256'h050505060606060707070708080808090909090A0A0A0B0B0B0B0C0C0C0C0D0D;
defparam prom_inst_2.INIT_RAM_35 = 256'hFCFDFDFDFDFEFEFEFEFFFFFFFF00000001010101020202020303030304040404;
defparam prom_inst_2.INIT_RAM_36 = 256'hF4F4F4F4F5F5F5F6F6F6F6F7F7F7F7F8F8F8F9F9F9F9FAFAFAFAFBFBFBFBFCFC;
defparam prom_inst_2.INIT_RAM_37 = 256'hEBEBEBECECECEDEDEDEDEEEEEEEEEFEFEFF0F0F0F0F1F1F1F1F2F2F2F3F3F3F3;
defparam prom_inst_2.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000E8E9E9E9E9EAEAEAEB;
defparam prom_inst_2.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[23:0],dout[31:24]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 8;
defparam prom_inst_3.RESET_MODE = "ASYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'h2F99046ED943AD1882EC56C02B95FF69D33DA7117BE54EB8228CF55FC9329C06;
defparam prom_inst_3.INIT_RAM_01 = 256'hCD38A4107BE752BD2994FF6BD641AC1782ED58C32E99046FDA44AF1A85EF5AC4;
defparam prom_inst_3.INIT_RAM_02 = 256'h44B11E8BF864D13EAA1783F05CC935A10E7AE652BE2A96026EDA46B21E8AF561;
defparam prom_inst_3.INIT_RAM_03 = 256'h90FF6DDB49B826940270DE4BB927950270DE4BB92694016EDC49B62390FD6AD7;
defparam prom_inst_3.INIT_RAM_04 = 256'hAD1D8DFC6CDC4BBB2A9A0979E857C736A51483F261D03FAD1C8BFA68D745B422;
defparam prom_inst_3.INIT_RAM_05 = 256'h950678E95BCC3DAF20910273E455C637A81889FA6ADB4BBC2C9C0C7DED5DCD3D;
defparam prom_inst_3.INIT_RAM_06 = 256'h43B72A9D1184F76ADD50C336A91C8E0173E658CB3DAF22940678EA5CCE40B123;
defparam prom_inst_3.INIT_RAM_07 = 256'hB4299F1489FF74E95ED348BD31A61B8F0478EC61D549BD31A5198D0175E95CD0;
defparam prom_inst_3.INIT_RAM_08 = 256'hE25AD149C037AF269D148B0279F066DD54CA41B72DA41A90067CF268DD53C93E;
defparam prom_inst_3.INIT_RAM_09 = 256'hC943BD36B02AA31D961089027BF46DE65FD750C941BA32AA239B138B037BF36A;
defparam prom_inst_3.INIT_RAM_0A = 256'h64E05DD955D14DC945C03CB733AE2AA5209B16910C87027CF772EC66E15BD54F;
defparam prom_inst_3.INIT_RAM_0B = 256'hAE2DAC2BA928A725A322A01E9C1A981693118F0C890784017EFB78F572EE6BE7;
defparam prom_inst_3.INIT_RAM_0C = 256'hA325A628A92BAC2DAE2FB031B232B333B434B434B434B434B433B332B231B02F;
defparam prom_inst_3.INIT_RAM_0D = 256'h3EC347CC50D458DC60E468EB6FF276F97CFF8205880B8E10931597199C1EA021;
defparam prom_inst_3.INIT_RAM_0E = 256'h7B028A119920A72EB53CC249CF56DC62E96FF57B00860C91169C21A62BB035BA;
defparam prom_inst_3.INIT_RAM_0F = 256'h54DF69F47E09931DA731BB45CE58E16BF47D068F18A129B23BC34BD35BE36BF3;
defparam prom_inst_3.INIT_RAM_10 = 256'hC553E16FFD8A18A533C04DDA67F4810D9A26B23FCB57E36EFA86119D28B33EC9;
defparam prom_inst_3.INIT_RAM_11 = 256'hCA5BED7E0FA031C253E474059525B545D565F58414A332C251E06EFD8C1AA937;
defparam prom_inst_3.INIT_RAM_12 = 256'h5DF2871CB146DA6F03972BBF53E77B0EA235C85BEE8114A739CC5EF08214A638;
defparam prom_inst_3.INIT_RAM_13 = 256'h7A13AC45DD760EA63ED66E069D35CC64FB9229BF56ED8319B046DC71079D32C8;
defparam prom_inst_3.INIT_RAM_14 = 256'h1DBA57F3902CC864009C38D36F0AA540DB7611AB46E07B15AF49E27C15AF48E1;
defparam prom_inst_3.INIT_RAM_15 = 256'h40E18223C36404A444E48323C26201A03FDE7C1BB958F69432D06D0BA946E380;
defparam prom_inst_3.INIT_RAM_16 = 256'hE0852ACF7318BC6105A94DF09437DB7E21C46709AC4EF19335D7791ABC5DFE9F;
defparam prom_inst_3.INIT_RAM_17 = 256'hF7A04AF39C45ED963EE78F37DF862ED67D24CB7219C0660DB359FFA54AF0963B;
defparam prom_inst_3.INIT_RAM_18 = 256'h812FDC8A37E5923FEC9945F29E4AF6A24EF9A550FBA751FCA751FCA650FAA44E;
defparam prom_inst_3.INIT_RAM_19 = 256'h792BDE9042F4A65709BA6B1CCD7E2FDF8F3FEF9F4FFFAE5D0DBC6B19C87625D3;
defparam prom_inst_3.INIT_RAM_1A = 256'hDA914900B66D24DA9046FCB2681DD2883DF1A65B0FC3782CDF9347FAAD6013C6;
defparam prom_inst_3.INIT_RAM_1B = 256'hA05D19D5904C07C37E39F3AE6923DD97510BC47E37F0A9621AD38B43FBB36B23;
defparam prom_inst_3.INIT_RAM_1C = 256'hC788490ACB8C4C0CCC8C4C0CCB8B4A09C8874504C2803EFCB97734F1AE6B28E4;
defparam prom_inst_3.INIT_RAM_1D = 256'h490FD69C6228EDB3783D02C78C5015D99D6124E8AB6E31F4B77A3CFEC0824405;
defparam prom_inst_3.INIT_RAM_1E = 256'h22EEB985501BE6B17C4611DBA56E3802CB945D26EEB77F470FD79F662DF4BB82;
defparam prom_inst_3.INIT_RAM_1F = 256'h4D1EF0C191623203D3A3734212E1B07F4E1CEAB9875522F0BD8A5724F1BD8A56;
defparam prom_inst_3.INIT_RAM_20 = 256'hC69D744B21F7CDA3794E24F9CEA3774C20F4C89C704316E9BC8F623406D8AA7C;
defparam prom_inst_3.INIT_RAM_21 = 256'h8865421EFAD6B28E69441FFAD5B08A643E18F2CBA57E572F08E0B991694018EF;
defparam prom_inst_3.INIT_RAM_22 = 256'h8F71543618FADCBE9F8061422303E3C3A38362422100DFBD9C7A583613F1CEAB;
defparam prom_inst_3.INIT_RAM_23 = 256'hD5BEA68F775F472E16FDE4CBB1987E644A3015FBE0C5AA8E72573B1E02E6C9AC;
defparam prom_inst_3.INIT_RAM_24 = 256'h5645342311FFEDDBC9B6A3907D6A56432F1A06F2DDC8B39D88725C46301A03EC;
defparam prom_inst_3.INIT_RAM_25 = 256'h0F04F9EEE3D7CCC0B4A79B8E8174675A4C3E30221305F6E7D8C8B8A999887867;
defparam prom_inst_3.INIT_RAM_26 = 256'hF9F5F0ECE7E2DDD7D2CCC6C0B9B3ACA59E968F877F776E655D544A41372D2319;
defparam prom_inst_3.INIT_RAM_27 = 256'h10131517191B1C1D1E1F2020202020201F1E1D1C1A19171512100D0A070400FD;
defparam prom_inst_3.INIT_RAM_28 = 256'h505A636C747D858D959CA4ABB2B9BFC5CCD1D7DDE2E7ECF0F5F9FD0104070B0D;
defparam prom_inst_3.INIT_RAM_29 = 256'hB5C5D5E5F5041322313F4D5B697784919EABB8C4D0DCE8F3FE09141F29333D47;
defparam prom_inst_3.INIT_RAM_2A = 256'h3950677E95ABC2D7ED03182D42576B7F93A7BBCEE1F407192B3D4F60728394A4;
defparam prom_inst_3.INIT_RAM_2B = 256'hD8F71533516E8CA9C6E3FF1B38536F8AA5C0DBF5102A435D768FA8C1D9F20A21;
defparam prom_inst_3.INIT_RAM_2C = 256'h8EB3D9FF24496E92B6DAFE2245688BAED0F2143658799ABBDBFC1C3C5C7B9AB9;
defparam prom_inst_3.INIT_RAM_2D = 256'h5582AFDC0936628EBAE5103B6691BBE50F39628BB4DD062E567EA5CCF41A4167;
defparam prom_inst_3.INIT_RAM_2E = 256'h295F93C8FC306498CBFE316496C9FB2C5E8FC0F1215282B1E1103F6E9DCBF927;
defparam prom_inst_3.INIT_RAM_2F = 256'h074480BDF93570ACE7225C97D10B457EB7F029619AD2094178AFE61C5389BFF4;
defparam prom_inst_3.INIT_RAM_30 = 256'hE82D72B6FA3E81C5084B8DCF115395D6175899D9195998D8175694D3114F8CCA;
defparam prom_inst_3.INIT_RAM_31 = 256'hC91663AFFB4793DE2974BF09539DE73079C20A539BE32A72B9FF468CD2185EA3;
defparam prom_inst_3.INIT_RAM_32 = 256'hA5FA4FA4F84CA0F4479AED3F92E43587D8297ACA1B6ABA0A59A8F64593E12F7C;
defparam prom_inst_3.INIT_RAM_33 = 256'h78D5328FEC48A5015CB8136EC8227DD63089E23B93EC449BF34AA1F84EA4FA50;
defparam prom_inst_3.INIT_RAM_34 = 256'h3CA2086DD2379C0064C82C8FF255B81A7CDE3FA00162C22282E241A0FF5EBC1A;
defparam prom_inst_3.INIT_RAM_35 = 256'hEE5CCB39A71482EF5BC834A00C77E24DB7228CF65FC8319A026BD23AA1086FD6;
defparam prom_inst_3.INIT_RAM_36 = 256'h880077EE64DB51C73CB1269B0F83F76BDE51C436A91B8CFE6FE050C030A0107F;
defparam prom_inst_3.INIT_RAM_37 = 256'h07870887078605840280FE7CF976F36FEB67E35ED954CF49C33CB62FA8209911;
defparam prom_inst_3.INIT_RAM_38 = 256'h000000000000000000000000000000000000000000000077FA7DFF8103840586;
defparam prom_inst_3.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_4 (
    .DO({prom_inst_4_dout_w[23:0],dout[39:32]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_4.READ_MODE = 1'b0;
defparam prom_inst_4.BIT_WIDTH = 8;
defparam prom_inst_4.RESET_MODE = "ASYNC";
defparam prom_inst_4.INIT_RAM_00 = 256'h69482807E6C6A58564432302E2C1A0805F3F1EFEDDBC9C7B5B3A19F9D8B89777;
defparam prom_inst_4.INIT_RAM_01 = 256'h7B5B3A1AF9D8B89777563515F4D4B39372513110F0CFAF8E6D4D2C0CEBCAAA89;
defparam prom_inst_4.INIT_RAM_02 = 256'h8E6D4D2C0BEBCAAA8969482707E6C6A58564432302E2C1A1805F3F1EFEDDBC9C;
defparam prom_inst_4.INIT_RAM_03 = 256'hA07F5F3E1EFDDDBC9C7B5A3A19F9D8B89776563515F4D4B39272513110EFCFAE;
defparam prom_inst_4.INIT_RAM_04 = 256'hB2927150300FEFCEAE8D6D4C2B0BEACAA98968472706E6C5A58463432202E1C1;
defparam prom_inst_4.INIT_RAM_05 = 256'hC4A48362422101E0C09F7F5E3D1DFCDCBB9B7A593918F8D7B79676553414F3D3;
defparam prom_inst_4.INIT_RAM_06 = 256'hD6B59574543312F2D1B190704F2F0EEECDAC8C6B4B2A0AE9C9A88767462605E5;
defparam prom_inst_4.INIT_RAM_07 = 256'hE7C7A68665442403E3C2A281614020FFDFBE9D7D5C3C1BFBDABA9979583717F6;
defparam prom_inst_4.INIT_RAM_08 = 256'hF8D8B79776563515F4D4B39372513110F0CFAF8E6E4D2D0CECCBAA8A69492808;
defparam prom_inst_4.INIT_RAM_09 = 256'h09E9C8A88767462605E5C4A48362422101E0C09F7F5E3E1DFDDCBC9B7B5A3919;
defparam prom_inst_4.INIT_RAM_0A = 256'h1AF9D9B89877573616F5D5B49473533212F1D1B0906F4F2E0DEDCCAC8B6B4A2A;
defparam prom_inst_4.INIT_RAM_0B = 256'h2A0AE9C9A88867472606E5C5A48463432202E1C1A0805F3F1EFDDDBC9C7B5B3A;
defparam prom_inst_4.INIT_RAM_0C = 256'h3A1AF9D9B89877573616F5D5B49473533212F1D1B0906F4F2E0EEDCDAC8C6B4B;
defparam prom_inst_4.INIT_RAM_0D = 256'h4A2909E8C8A78766462505E4C4A38362422101E1C0A07F5F3E1EFDDDBC9C7B5B;
defparam prom_inst_4.INIT_RAM_0E = 256'h593918F8D7B79676553514F4D3B39272513110F0D0AF8F6E4E2D0DECCCAB8B6A;
defparam prom_inst_4.INIT_RAM_0F = 256'h68472706E6C6A58564442303E2C2A181604020FFDFBE9E7D5D3C1CFBDBBA9A79;
defparam prom_inst_4.INIT_RAM_10 = 256'h76563515F4D4B49373523211F1D0B0906F4F2E0EEDCDAC8C6B4B2B0AEAC9A988;
defparam prom_inst_4.INIT_RAM_11 = 256'h8464432303E2C2A181604020FFDFBE9E7D5D3C1CFCDBBB9A7A593918F8D8B797;
defparam prom_inst_4.INIT_RAM_12 = 256'h9271513110F0CFAF8F6E4E2D0DECCCAC8B6B4A2A09E9C9A88867472606E6C5A5;
defparam prom_inst_4.INIT_RAM_13 = 256'h9F7F5E3E1DFDDDBC9C7B5B3B1AFAD9B99878583717F6D6B69575543414F3D3B2;
defparam prom_inst_4.INIT_RAM_14 = 256'hAC8B6B4A2A0AE9C9A98868472707E6C6A58565442403E3C3A28261412100E0BF;
defparam prom_inst_4.INIT_RAM_15 = 256'hB89777573616F6D5B59474543313F3D2B29171513010EFCFAF8E6E4E2D0DECCC;
defparam prom_inst_4.INIT_RAM_16 = 256'hC3A38362422201E1C1A0805F3F1FFEDEBE9D7D5D3C1CFBDBBB9A7A5A3919F8D8;
defparam prom_inst_4.INIT_RAM_17 = 256'hCEAE8E6D4D2D0CECCCAB8B6B4A2A0AE9C9A98868482707E7C6A68565452404E4;
defparam prom_inst_4.INIT_RAM_18 = 256'hD9B99878583717F7D6B69675553514F4D4B39373523212F1D1B19070502F0FEF;
defparam prom_inst_4.INIT_RAM_19 = 256'hE3C3A28262412101E1C0A0805F3F1FFEDEBE9D7D5D3C1CFCDCBB9B7B5A3A1AF9;
defparam prom_inst_4.INIT_RAM_1A = 256'hECCCAC8C6B4B2B0AEACAA98969492808E8C7A78767462606E5C5A58464442403;
defparam prom_inst_4.INIT_RAM_1B = 256'hF5D5B59474543413F3D3B29272523111F1D1B090704F2F0FEFCEAE8E6D4D2D0D;
defparam prom_inst_4.INIT_RAM_1C = 256'hFDDDBD9D7C5C3C1CFBDBBB9B7A5A3A1AF9D9B99978583817F7D7B79676563615;
defparam prom_inst_4.INIT_RAM_1D = 256'h05E5C4A48464432303E3C3A28262422101E1C1A08060401FFFDFBF9E7E5E3E1E;
defparam prom_inst_4.INIT_RAM_1E = 256'h0CEBCBAB8B6B4A2A0AEACAA98969492908E8C8A88767472707E6C6A686654525;
defparam prom_inst_4.INIT_RAM_1F = 256'h12F2D1B19171513110F0D0B0906F4F2F0FEFCEAE8E6E4E2D0DEDCDAD8C6C4C2C;
defparam prom_inst_4.INIT_RAM_20 = 256'h17F7D7B79776563616F6D6B59575553515F4D4B49474543313F3D3B393725232;
defparam prom_inst_4.INIT_RAM_21 = 256'h1CFCDCBC9B7B5B3B1BFBDBBA9A7A5A3A1AFAD9B99979593919F8D8B898785837;
defparam prom_inst_4.INIT_RAM_22 = 256'h2000E0C0A07F5F3F1FFFDFBF9F7F5E3E1EFEDEBE9E7E5D3D1DFDDDBD9D7C5C3C;
defparam prom_inst_4.INIT_RAM_23 = 256'h2303E3C3A38363432302E2C2A28262422202E2C1A18161412101E1C1A1806040;
defparam prom_inst_4.INIT_RAM_24 = 256'h2606E6C6A68565452505E5C5A58565452505E5C4A48464442404E4C4A4846443;
defparam prom_inst_4.INIT_RAM_25 = 256'h2808E7C7A78767472707E7C7A78767472707E7C7A78766462606E6C6A6866646;
defparam prom_inst_4.INIT_RAM_26 = 256'h2808E8C8A88868482808E8C8A88868482808E8C8A88868482808E8C8A8886848;
defparam prom_inst_4.INIT_RAM_27 = 256'h2909E9C9A98969492909E9C9A98969492909E9C9A98969492909E9C9A9896948;
defparam prom_inst_4.INIT_RAM_28 = 256'h2808E8C8A88868482808E8C8A88868482808E8C8A88868482808E8C9A9896949;
defparam prom_inst_4.INIT_RAM_29 = 256'h2606E6C6A68767472707E7C7A78767472707E7C7A78767472708E8C8A8886848;
defparam prom_inst_4.INIT_RAM_2A = 256'h2404E4C4A48464442405E5C5A58565452505E5C5A58566462606E6C6A6866646;
defparam prom_inst_4.INIT_RAM_2B = 256'h2000E1C1A18161412101E1C2A28262422202E2C2A38363432303E3C3A3836444;
defparam prom_inst_4.INIT_RAM_2C = 256'h1CFCDCBC9D7D5D3D1DFDDDBE9E7E5E3E1EFEDFBF9F7F5F3F1FFFE0C0A0806040;
defparam prom_inst_4.INIT_RAM_2D = 256'h17F7D7B79878583818F8D9B9997959391AFADABA9A7A5B3B1BFBDBBB9B7C5C3C;
defparam prom_inst_4.INIT_RAM_2E = 256'h11F1D1B19172523212F2D3B39373533414F4D4B49575553515F6D6B696765637;
defparam prom_inst_4.INIT_RAM_2F = 256'h0AEACAAA8A6B4B2B0BECCCAC8C6D4D2D0DEDCEAE8E6E4F2F0FEFCFB090705030;
defparam prom_inst_4.INIT_RAM_30 = 256'h01E2C2A28263432304E4C4A48565452506E6C6A68767472708E8C8A889694929;
defparam prom_inst_4.INIT_RAM_31 = 256'hF8D9B999795A3A1AFBDBBB9C7C5C3C1DFDDDBE9E7E5E3F1FFFDFC0A080614121;
defparam prom_inst_4.INIT_RAM_32 = 256'hEECEAF8F6F503010F1D1B19272523313F3D4B49475553516F6D6B69777573818;
defparam prom_inst_4.INIT_RAM_33 = 256'hE3C3A48464452506E6C6A78767482808E9C9A98A6A4A2B0BEBCCAC8C6D4D2D0E;
defparam prom_inst_4.INIT_RAM_34 = 256'hD7B79878583919FADABA9B7B5B3C1CFDDDBD9E7E5F3F1F00E0C0A18161422203;
defparam prom_inst_4.INIT_RAM_35 = 256'hC9AA8A6B4B2C0CECCDAD8E6E4F2F0FF0D0B19171523213F3D4B49475553616F6;
defparam prom_inst_4.INIT_RAM_36 = 256'hBB9C7C5C3D1DFEDEBF9F8060412101E2C2A38364442505E5C6A68767482809E9;
defparam prom_inst_4.INIT_RAM_37 = 256'hAC8C6D4D2E0EEFCFB09070513112F2D3B39474553516F6D7B7987859391AFADB;
defparam prom_inst_4.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000C7A78868492A0AEBCB;
defparam prom_inst_4.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_5 (
    .DO({prom_inst_5_dout_w[23:0],dout[47:40]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_5.READ_MODE = 1'b0;
defparam prom_inst_5.BIT_WIDTH = 8;
defparam prom_inst_5.RESET_MODE = "ASYNC";
defparam prom_inst_5.INIT_RAM_00 = 256'h1D1D1D1D1C1C1C1C1C1C1C1C1B1B1B1B1B1B1B1A1A1A1A1A1A1A1A1919191919;
defparam prom_inst_5.INIT_RAM_01 = 256'h2121212120202020202020201F1F1F1F1F1F1F1F1E1E1E1E1E1E1E1E1D1D1D1D;
defparam prom_inst_5.INIT_RAM_02 = 256'h2525252525242424242424242423232323232323232222222222222221212121;
defparam prom_inst_5.INIT_RAM_03 = 256'h2929292929282828282828282827272727272727272626262626262626252525;
defparam prom_inst_5.INIT_RAM_04 = 256'h2D2D2D2D2D2D2C2C2C2C2C2C2C2C2B2B2B2B2B2B2B2B2A2A2A2A2A2A2A2A2929;
defparam prom_inst_5.INIT_RAM_05 = 256'h31313131313131303030303030302F2F2F2F2F2F2F2F2E2E2E2E2E2E2E2E2D2D;
defparam prom_inst_5.INIT_RAM_06 = 256'h3535353535353534343434343434343333333333333333323232323232323231;
defparam prom_inst_5.INIT_RAM_07 = 256'h3939393939393939383838383838383737373737373737363636363636363635;
defparam prom_inst_5.INIT_RAM_08 = 256'h3D3D3D3D3D3D3D3D3C3C3C3C3C3C3C3C3B3B3B3B3B3B3B3B3A3A3A3A3A3A3A3A;
defparam prom_inst_5.INIT_RAM_09 = 256'h42414141414141414140404040404040403F3F3F3F3F3F3F3E3E3E3E3E3E3E3E;
defparam prom_inst_5.INIT_RAM_0A = 256'h4645454545454545454444444444444444434343434343434342424242424242;
defparam prom_inst_5.INIT_RAM_0B = 256'h4A4A494949494949494948484848484848484747474747474746464646464646;
defparam prom_inst_5.INIT_RAM_0C = 256'h4E4E4D4D4D4D4D4D4D4D4C4C4C4C4C4C4C4C4B4B4B4B4B4B4B4B4A4A4A4A4A4A;
defparam prom_inst_5.INIT_RAM_0D = 256'h525252515151515151515150505050505050504F4F4F4F4F4F4F4E4E4E4E4E4E;
defparam prom_inst_5.INIT_RAM_0E = 256'h5656565555555555555555545454545454545453535353535353535252525252;
defparam prom_inst_5.INIT_RAM_0F = 256'h5A5A5A5A59595959595959595858585858585857575757575757575656565656;
defparam prom_inst_5.INIT_RAM_10 = 256'h5E5E5E5E5D5D5D5D5D5D5D5D5C5C5C5C5C5C5C5C5B5B5B5B5B5B5B5B5A5A5A5A;
defparam prom_inst_5.INIT_RAM_11 = 256'h62626262626161616161616160606060606060605F5F5F5F5F5F5F5F5E5E5E5E;
defparam prom_inst_5.INIT_RAM_12 = 256'h6666666666656565656565656564646464646464646363636363636363626262;
defparam prom_inst_5.INIT_RAM_13 = 256'h6A6A6A6A6A696969696969696968686868686868686767676767676767666666;
defparam prom_inst_5.INIT_RAM_14 = 256'h6E6E6E6E6E6E6D6D6D6D6D6D6D6D6C6C6C6C6C6C6C6C6B6B6B6B6B6B6B6B6A6A;
defparam prom_inst_5.INIT_RAM_15 = 256'h727272727272717171717171717170707070707070706F6F6F6F6F6F6F6F6E6E;
defparam prom_inst_5.INIT_RAM_16 = 256'h7676767676767675757575757575747474747474747473737373737373737272;
defparam prom_inst_5.INIT_RAM_17 = 256'h7A7A7A7A7A7A7A79797979797979797878787878787878777777777777777776;
defparam prom_inst_5.INIT_RAM_18 = 256'h7E7E7E7E7E7E7E7D7D7D7D7D7D7D7D7C7C7C7C7C7C7C7C7B7B7B7B7B7B7B7B7A;
defparam prom_inst_5.INIT_RAM_19 = 256'h82828282828282828181818181818180808080808080807F7F7F7F7F7F7F7F7E;
defparam prom_inst_5.INIT_RAM_1A = 256'h8686868686868686858585858585858584848484848484848383838383838383;
defparam prom_inst_5.INIT_RAM_1B = 256'h8A8A8A8A8A8A8A8A898989898989898988888888888888888787878787878787;
defparam prom_inst_5.INIT_RAM_1C = 256'h8E8E8E8E8E8E8E8E8D8D8D8D8D8D8D8D8C8C8C8C8C8C8C8C8B8B8B8B8B8B8B8B;
defparam prom_inst_5.INIT_RAM_1D = 256'h9392929292929292929191919191919191909090909090908F8F8F8F8F8F8F8F;
defparam prom_inst_5.INIT_RAM_1E = 256'h9796969696969696969595959595959595949494949494949493939393939393;
defparam prom_inst_5.INIT_RAM_1F = 256'h9B9A9A9A9A9A9A9A9A9999999999999999989898989898989897979797979797;
defparam prom_inst_5.INIT_RAM_20 = 256'h9F9E9E9E9E9E9E9E9E9D9D9D9D9D9D9D9D9C9C9C9C9C9C9C9C9B9B9B9B9B9B9B;
defparam prom_inst_5.INIT_RAM_21 = 256'hA3A2A2A2A2A2A2A2A2A1A1A1A1A1A1A1A1A0A0A0A0A0A0A0A09F9F9F9F9F9F9F;
defparam prom_inst_5.INIT_RAM_22 = 256'hA7A7A6A6A6A6A6A6A6A5A5A5A5A5A5A5A5A4A4A4A4A4A4A4A4A3A3A3A3A3A3A3;
defparam prom_inst_5.INIT_RAM_23 = 256'hABABAAAAAAAAAAAAAAAAA9A9A9A9A9A9A9A9A8A8A8A8A8A8A8A8A7A7A7A7A7A7;
defparam prom_inst_5.INIT_RAM_24 = 256'hAFAFAEAEAEAEAEAEAEAEADADADADADADADADACACACACACACACACABABABABABAB;
defparam prom_inst_5.INIT_RAM_25 = 256'hB3B3B2B2B2B2B2B2B2B2B1B1B1B1B1B1B1B1B0B0B0B0B0B0B0B0AFAFAFAFAFAF;
defparam prom_inst_5.INIT_RAM_26 = 256'hB7B7B6B6B6B6B6B6B6B6B5B5B5B5B5B5B5B5B4B4B4B4B4B4B4B4B3B3B3B3B3B3;
defparam prom_inst_5.INIT_RAM_27 = 256'hBBBBBABABABABABABABAB9B9B9B9B9B9B9B9B8B8B8B8B8B8B8B8B7B7B7B7B7B7;
defparam prom_inst_5.INIT_RAM_28 = 256'hBFBFBEBEBEBEBEBEBEBEBDBDBDBDBDBDBDBDBCBCBCBCBCBCBCBCBBBBBBBBBBBB;
defparam prom_inst_5.INIT_RAM_29 = 256'hC3C3C2C2C2C2C2C2C2C2C1C1C1C1C1C1C1C1C0C0C0C0C0C0C0C0BFBFBFBFBFBF;
defparam prom_inst_5.INIT_RAM_2A = 256'hC7C7C6C6C6C6C6C6C6C6C5C5C5C5C5C5C5C5C4C4C4C4C4C4C4C4C3C3C3C3C3C3;
defparam prom_inst_5.INIT_RAM_2B = 256'hCBCBCACACACACACACACAC9C9C9C9C9C9C9C9C8C8C8C8C8C8C8C8C7C7C7C7C7C7;
defparam prom_inst_5.INIT_RAM_2C = 256'hCFCECECECECECECECECDCDCDCDCDCDCDCDCCCCCCCCCCCCCCCCCBCBCBCBCBCBCB;
defparam prom_inst_5.INIT_RAM_2D = 256'hD3D2D2D2D2D2D2D2D2D1D1D1D1D1D1D1D1D0D0D0D0D0D0D0D0CFCFCFCFCFCFCF;
defparam prom_inst_5.INIT_RAM_2E = 256'hD7D6D6D6D6D6D6D6D6D5D5D5D5D5D5D5D5D4D4D4D4D4D4D4D4D3D3D3D3D3D3D3;
defparam prom_inst_5.INIT_RAM_2F = 256'hDBDADADADADADADADAD9D9D9D9D9D9D9D9D8D8D8D8D8D8D8D8D7D7D7D7D7D7D7;
defparam prom_inst_5.INIT_RAM_30 = 256'hDFDEDEDEDEDEDEDEDEDDDDDDDDDDDDDDDDDCDCDCDCDCDCDCDCDBDBDBDBDBDBDB;
defparam prom_inst_5.INIT_RAM_31 = 256'hE2E2E2E2E2E2E2E2E1E1E1E1E1E1E1E1E0E0E0E0E0E0E0E0DFDFDFDFDFDFDFDF;
defparam prom_inst_5.INIT_RAM_32 = 256'hE6E6E6E6E6E6E6E6E5E5E5E5E5E5E5E5E4E4E4E4E4E4E4E4E3E3E3E3E3E3E3E3;
defparam prom_inst_5.INIT_RAM_33 = 256'hEAEAEAEAEAEAEAEAE9E9E9E9E9E9E9E9E8E8E8E8E8E8E8E8E7E7E7E7E7E7E7E7;
defparam prom_inst_5.INIT_RAM_34 = 256'hEEEEEEEEEEEEEEEDEDEDEDEDEDEDEDECECECECECECECECECEBEBEBEBEBEBEBEB;
defparam prom_inst_5.INIT_RAM_35 = 256'hF2F2F2F2F2F2F2F1F1F1F1F1F1F1F1F0F0F0F0F0F0F0F0EFEFEFEFEFEFEFEFEE;
defparam prom_inst_5.INIT_RAM_36 = 256'hF6F6F6F6F6F6F5F5F5F5F5F5F5F5F5F4F4F4F4F4F4F4F4F3F3F3F3F3F3F3F3F2;
defparam prom_inst_5.INIT_RAM_37 = 256'hFAFAFAFAFAFAF9F9F9F9F9F9F9F9F8F8F8F8F8F8F8F8F7F7F7F7F7F7F7F7F6F6;
defparam prom_inst_5.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000FBFBFBFBFBFBFBFAFA;
defparam prom_inst_5.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule //coef_prom
